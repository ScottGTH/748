import uvm_pkg::*;
`include "uvm_macros.svh"

import decode_in_pkg::*;
import decode_out_pkg::*;
import decode_test_pkg::*;

module hvl_top();

    initial run_test();
endmodule