package decode_out_pkg;
   
   import uvm_pkg::*;
   import para_type_pkg::*;

   `include "uvm_macros.svh"

   `include "src/decode_out_transaction.svh"

   `include "src/decode_out_configuration.svh"
   `include "src/decode_out_monitor.svh"

   `include "src/decode_out_transaction_coverage.svh"
   `include "src/decode_out_agent.svh"

endpackage

